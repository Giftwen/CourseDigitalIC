/*
 * @Author: WenJiaBao-2022E8020282071
 * @Date: 2022-10-12 23:40:14
 * @LastEditTime: 2022-10-12 23:42:01
 * @Description: 
 * 
 * Copyright (c) 2022 by WenJiaBao wenjiabao0919@163.com, All Rights Reserved. 
 */
 module watch(
    input
 );
