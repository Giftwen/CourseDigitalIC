/*
 * @Author: WenJiaBao-2022E8020282071
 * @Date: 2022-10-18 17:21:22
 * @LastEditTime: 2022-10-18 17:28:18
 * @Description: 
 * 
 * Copyright (c) 2022 by WenJiaBao wenjiabao0919@163.com, All Rights Reserved. 
 */
module barrel(
    input   [15:0]  a_i,
    input   [15:0]  b_i,
    output  [16:0]  sum_o
);

endmodule