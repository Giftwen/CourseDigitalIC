module decode16_5(
    input       [4:0]   in   ,
    output reg [15:0]   out
);

always @(*) begin
    case(in)
        5'b00000:out<=16'b0000_0000_0000_0000;
        5'b00001:out<=16'b0000_0000_0000_0001;
        5'b00010:out<=16'b0000_0000_0000_0011;
        5'b00011:out<=16'b0000_0000_0000_0111;
        5'b00100:out<=16'b0000_0000_0000_1111;
        5'b00101:out<=16'b0000_0000_0001_1111;
        5'b00110:out<=16'b0000_0000_0011_1111;
        5'b00111:out<=16'b0000_0000_0111_1111;
        5'b01000:out<=16'b0000_0000_1111_1111;
        5'b01001:out<=16'b0000_0001_1111_1111;
        5'b01010:out<=16'b0000_0011_1111_1111;
        5'b01011:out<=16'b0000_0111_1111_1111;
        5'b01100:out<=16'b0000_1111_1111_1111;
        5'b01101:out<=16'b0001_1111_1111_1111;
        5'b01110:out<=16'b0011_1111_1111_1111;
        5'b01111:out<=16'b0111_1111_1111_1111;
        5'b10000:out<=16'b1111_1111_1111_1111;
        default:begin
            out<=16'b0000_0000_0000;
        end
    endcase
end

endmodule