/*
 * @Author: WenJiaBao-2022E8020282071
 * @Date: 2022-10-12 23:40:02
 * @LastEditTime: 2022-10-12 23:41:49
 * @Description: 
 * 
 * Copyright (c) 2022 by WenJiaBao wenjiabao0919@163.com, All Rights Reserved. 
 */
 module clk_gen();
